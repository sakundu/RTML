`define INPUT_BITWIDTH xx_ip_bitwidth_xx
`define BITWIDTH xx_bitwidth_xx
`define NUM_CYCLE xx_num_cycle_xx
`define LOG_NUM_CYCLE xx_log_num_cycle_xx
`define SIZE xx_size_xx
`define NUMBER_UNIT xx_unit_xx
`define INST_BITWIDTH 4

// `define SVM 1
// `define LINEAR 1
// `define LOGISTIC 1
// `define RECO 1
